module deserializer (CLK , RST , sampled_bit , deser_en  , P_DATA);

////////////////////////////////////////////////////////
/////////////////// IN/OUT PORTS /////////////////////// 
////////////////////////////////////////////////////////

input							CLK;
input							RST;
input							sampled_bit;
input							deser_en;
output reg 		[63:0] 			P_DATA;

////////////////////////////////////////////////////////
///////////////// Internal signals ///////////////////// 
////////////////////////////////////////////////////////

reg				[5:0] 			counter;
reg				[2:0]			index;
wire			[4:0]			sample_time;

////////////////////////////////////////////////////////
////////////////// ASSIGN STATMENTS //////////////////// 
////////////////////////////////////////////////////////

assign sample_time = 64;

////////////////////////////////////////////////////////
////////////////// Deserializing /////////////////////// 
////////////////////////////////////////////////////////

always @ (posedge CLK or negedge RST) begin
	if (!RST) begin
		P_DATA  <= 0;
		counter <= 0;
		index   <= 0;
	end
	else begin
		if (deser_en) begin
			if (counter != sample_time) begin
				P_DATA [index] <= sampled_bit;
				index <= index + 1;
			end
			counter <= counter + 1;
			if (counter == 64)
			counter <= 0;
		end
	end
end
endmodule 
